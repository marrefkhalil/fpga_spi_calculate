module spi_slave (


);